package seq_mult_pkg;

localparam DW       = 8;

endpackage: seq_mult_pkg
