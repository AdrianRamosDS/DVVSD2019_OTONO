package mdr_pkg;

localparam DW       	= 16;
localparam DW_DBL 	= 32;
localparam SQRT_NBitsForCounter = 5;

endpackage
